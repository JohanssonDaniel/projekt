library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.numeric_std.ALL;
--use ieee.numeric_bit;
--use ieee.numeric_std;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity myPC is
	port(
		clk,rst : in STD_LOGIC;
		k1,k2 : in STD_LOGIC_VECTOR(7 downto 0);
		SEQ : in STD_LOGIC_VECTOR(3 downto 0);
		my_out : out STD_LOGIC_VECTOR(7 downto 0)
	);
end myPC;

architecture Behavorial of myPC is 
	SIGNAL myCounter : STD_LOGIC_VECTOR(7 downto 0);
begin
	process(clk,rst) begin
		if rst = '1' then
				myCounter <= X"00";
		else
			case SEQ is
				when "0000" => myCounter <= myCounter + 1; 
				when "0001" => myCounter <= k1;
				when "0010" => myCounter <= k2;
				when "0011" => myCounter <= X"00";
				when others => myCounter <= myCounter;
			end case;
		end if;
	end process;
	
	my_out <= myCounter;
end Behavorial;
	
