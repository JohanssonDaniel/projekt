entity mymem is
 port(instructionset: out mymem);
end mymem;

architecture set of mymem is

begin  -- set

 type mymem is array (0 to 127) of std_logic_vector(27 downto 0);
 signal instructionset : mymem := (X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000",
                                   X"0000000");


end set;
